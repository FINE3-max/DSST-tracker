parameter IMG_width = 640;
parameter IMG_height = 480;

parameter Kuang_width = 300;
parameter Kuang_height = 150;

parameter Kuang_mid_x = 150;
parameter Kuang_mid_y = 75;

parameter Kuang_x_end = 490;//1280-150=1130//640-150=490
parameter Kuang_y_end = 405;//720-75=645//480-75=405